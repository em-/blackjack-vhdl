package vectors is
    type natural_vector is array(natural range <>) of natural;
    type boolean_vector is array(natural range <>) of boolean;
end vectors;
